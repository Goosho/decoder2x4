library verilog;
use verilog.vl_types.all;
entity decoder2x4_vlg_vec_tst is
end decoder2x4_vlg_vec_tst;
